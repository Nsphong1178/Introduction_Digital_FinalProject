entity HelloWorld is
end entity;

architecture lab of HelloWorld is
begin 

	process is
	begin 
		report "Hello Aloo";
		wait;
	end process;

end architecture;
